module instruction_decode_stage ();

endmodule
