package common_instructions_pkg;

  typedef enum logic [31:0] {
    // instr      =     func7____rs2___rs1_func3_rd___op_code,
    INSTR_LUI     = 32'b???????_?????_?????_???_?????_0110111,
    INSTR_AUIPC   = 32'b???????_?????_?????_???_?????_0010111,
    INSTR_JAL     = 32'b???????_?????_?????_???_?????_1101111,
    INSTR_JALR    = 32'b???????_?????_?????_000_?????_1100111,
    INSTR_BEQ     = 32'b???????_?????_?????_000_?????_1100011,
    INSTR_BNE     = 32'b???????_?????_?????_001_?????_1100011,
    INSTR_BLT     = 32'b???????_?????_?????_100_?????_1100011,
    INSTR_BGE     = 32'b???????_?????_?????_101_?????_1100011,
    INSTR_BLTU    = 32'b???????_?????_?????_110_?????_1100011,
    INSTR_BGEU    = 32'b???????_?????_?????_111_?????_1100011,
    INSTR_LB      = 32'b???????_?????_?????_000_?????_0000011,
    INSTR_LH      = 32'b???????_?????_?????_001_?????_0000011,
    INSTR_LW      = 32'b???????_?????_?????_010_?????_0000011,
    INSTR_LBU     = 32'b???????_?????_?????_100_?????_0000011,
    INSTR_LHU     = 32'b???????_?????_?????_101_?????_0000011,
    INSTR_SB      = 32'b???????_?????_?????_000_?????_0100011,
    INSTR_SH      = 32'b???????_?????_?????_001_?????_0100011,
    INSTR_SW      = 32'b???????_?????_?????_010_?????_0100011,
    INSTR_ADDI    = 32'b???????_?????_?????_000_?????_0010011,
    INSTR_SLTI    = 32'b???????_?????_?????_010_?????_0010011,
    INSTR_SLTIU   = 32'b???????_?????_?????_011_?????_0010011,
    INSTR_XORI    = 32'b???????_?????_?????_100_?????_0010011,
    INSTR_ORI     = 32'b???????_?????_?????_110_?????_0010011,
    INSTR_ANDI    = 32'b???????_?????_?????_111_?????_0010011,
    INSTR_SLLI    = 32'b0000000_?????_?????_001_?????_0010011,
    INSTR_SRLI    = 32'b0000000_?????_?????_101_?????_0010011,
    INSTR_SRAI    = 32'b0100000_?????_?????_101_?????_0010011,
    INSTR_ADD     = 32'b0000000_?????_?????_000_?????_0110011,
    INSTR_SUB     = 32'b0100000_?????_?????_000_?????_0110011,
    INSTR_SLL     = 32'b0000000_?????_?????_001_?????_0110011,
    INSTR_SLT     = 32'b0000000_?????_?????_010_?????_0110011,
    INSTR_SLTU    = 32'b0000000_?????_?????_011_?????_0110011,
    INSTR_XOR     = 32'b0000000_?????_?????_100_?????_0110011,
    INSTR_SRL     = 32'b0000000_?????_?????_101_?????_0110011,
    INSTR_SRA     = 32'b0100000_?????_?????_101_?????_0110011,
    INSTR_OR      = 32'b0000000_?????_?????_110_?????_0110011,
    INSTR_AND     = 32'b0000000_?????_?????_111_?????_0110011,
    INSTR_MUL     = 32'b0000001_?????_?????_000_?????_0110011,
    INSTR_MULH    = 32'b0000001_?????_?????_001_?????_0110011,
    INSTR_DIV     = 32'b0000001_?????_?????_100_?????_0110011,
    INSTR_DIVU    = 32'b0000001_?????_?????_101_?????_0110011,
    INSTR_REM     = 32'b0000001_?????_?????_110_?????_0110011,
    INSTR_REMU    = 32'b0000001_?????_?????_111_?????_0110011,
    INSTR_FLW     = 32'b???????_?????_?????_010_?????_0000111,
    INSTR_FSW     = 32'b???????_?????_?????_010_?????_0100111,
    INSTR_FADD_S  = 32'b0000000_?????_?????_???_?????_1010011,
    INSTR_FSUB_S  = 32'b0000100_?????_?????_???_?????_1010011,
    INSTR_FMUL_S  = 32'b0001000_?????_?????_???_?????_1010011,
    INSTR_FDIV_S  = 32'b0001100_?????_?????_???_?????_1010011,
    INSTR_FSQRT_S = 32'b0101100_00000_?????_???_?????_1010011,
    INSTR_FMV_X_W = 32'b1110000_00000_?????_000_?????_1010011,
    INSTR_FEQ_S   = 32'b1010000_?????_?????_010_?????_1010011,
    INSTR_FLT_S   = 32'b1010000_?????_?????_001_?????_1010011,
    INSTR_FLE_S   = 32'b1010000_?????_?????_000_?????_1010011,
    INSTR_FMV_W_X = 32'b1111000_00000_?????_000_?????_1010011,
    INSTR_HALT    = 32'b1111111_11111_11111_111_11111_1111111
  } normal_instructions_t;

  typedef enum logic [15:0] {
    INSTR_C_NOP  = 16'b000_0_00000_00000_01,
    INSTR_C_ADDI = 16'b000_?_?????_?????_01
  } compressed_instructions_t;

endpackage


