module writeback_stage ();

endmodule
