module memory_stage ();

endmodule
