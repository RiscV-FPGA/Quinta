`timescale 1ns / 1ps

module tb_top;

  logic clk = 0;
  logic rst = 1;

  integer cycle = 0;
  int test_length = 500;
  int clk_period = 10;

  top top_uut (
      .clk(clk),
      .rst(rst)
  );

  always #(clk_period / 2) clk = ~clk;
  always #clk_period cycle++;

  initial begin

    #(clk_period * 2);
    rst <= 0;

  end

  initial begin
    $dumpfile("waveform.vcd");
    $dumpvars(0, tb_top);
    $display("Done!");

    #test_length;  //test length

    $finish();
  end

endmodule
