module execute_stage ();

endmodule
