module instruction_fetch_stage ();

endmodule
